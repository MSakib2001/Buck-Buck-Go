// VGA.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module VGA (
		input  wire  clk_clk,                        //                      clk.clk
		input  wire  reset_reset_n,                  //                    reset.reset_n
		output wire  video_pll_0_reset_source_reset, // video_pll_0_reset_source.reset
		output wire  video_pll_0_vga_clk_clk         //      video_pll_0_vga_clk.clk
	);

	VGA_video_pll_0 video_pll_0 (
		.ref_clk_clk        (clk_clk),                        //      ref_clk.clk
		.ref_reset_reset    (~reset_reset_n),                 //    ref_reset.reset
		.vga_clk_clk        (video_pll_0_vga_clk_clk),        //      vga_clk.clk
		.reset_source_reset (video_pll_0_reset_source_reset)  // reset_source.reset
	);

endmodule
