
module VGA (
	clk_clk,
	reset_reset_n,
	video_pll_0_vga_clk_clk,
	video_pll_0_reset_source_reset);	

	input		clk_clk;
	input		reset_reset_n;
	output		video_pll_0_vga_clk_clk;
	output		video_pll_0_reset_source_reset;
endmodule
