// data_mem_2.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module data_mem_2 (
		input  wire        palette_clk1_clk,         //   palette_clk1.clk
		input  wire        palette_reset1_reset,     // palette_reset1.reset
		input  wire        palette_reset1_reset_req, //               .reset_req
		input  wire [5:0]  palette_s1_address,       //     palette_s1.address
		input  wire        palette_s1_clken,         //               .clken
		input  wire        palette_s1_chipselect,    //               .chipselect
		input  wire        palette_s1_write,         //               .write
		output wire [31:0] palette_s1_readdata,      //               .readdata
		input  wire [31:0] palette_s1_writedata,     //               .writedata
		input  wire [3:0]  palette_s1_byteenable     //               .byteenable
	);

	data_mem_2_palette palette (
		.clk        (palette_clk1_clk),         //   clk1.clk
		.address    (palette_s1_address),       //     s1.address
		.clken      (palette_s1_clken),         //       .clken
		.chipselect (palette_s1_chipselect),    //       .chipselect
		.write      (palette_s1_write),         //       .write
		.readdata   (palette_s1_readdata),      //       .readdata
		.writedata  (palette_s1_writedata),     //       .writedata
		.byteenable (palette_s1_byteenable),    //       .byteenable
		.reset      (palette_reset1_reset),     // reset1.reset
		.reset_req  (palette_reset1_reset_req), //       .reset_req
		.freeze     (1'b0)                      // (terminated)
	);

endmodule
