// RAM.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module RAM (
		input  wire        clk_ram_clk,          //   clk_ram.clk
		input  wire [9:0]  ram_slave_address,    // ram_slave.address
		input  wire        ram_slave_clken,      //          .clken
		input  wire        ram_slave_chipselect, //          .chipselect
		input  wire        ram_slave_write,      //          .write
		output wire [31:0] ram_slave_readdata,   //          .readdata
		input  wire [31:0] ram_slave_writedata,  //          .writedata
		input  wire [3:0]  ram_slave_byteenable, //          .byteenable
		input  wire        rst_ram_reset,        //   rst_ram.reset
		input  wire        rst_ram_reset_req     //          .reset_req
	);

	RAM_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_ram_clk),          //   clk1.clk
		.address    (ram_slave_address),    //     s1.address
		.clken      (ram_slave_clken),      //       .clken
		.chipselect (ram_slave_chipselect), //       .chipselect
		.write      (ram_slave_write),      //       .write
		.readdata   (ram_slave_readdata),   //       .readdata
		.writedata  (ram_slave_writedata),  //       .writedata
		.byteenable (ram_slave_byteenable), //       .byteenable
		.reset      (rst_ram_reset),        // reset1.reset
		.reset_req  (rst_ram_reset_req),    //       .reset_req
		.freeze     (1'b0)                  // (terminated)
	);

endmodule
