// background_data.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module background_data (
		input  wire        onchip_memory2_0_clk1_clk,         //   onchip_memory2_0_clk1.clk
		input  wire        onchip_memory2_0_reset1_reset,     // onchip_memory2_0_reset1.reset
		input  wire        onchip_memory2_0_reset1_reset_req, //                        .reset_req
		input  wire [18:0] onchip_memory2_0_s1_address,       //     onchip_memory2_0_s1.address
		input  wire        onchip_memory2_0_s1_debugaccess,   //                        .debugaccess
		input  wire        onchip_memory2_0_s1_clken,         //                        .clken
		input  wire        onchip_memory2_0_s1_chipselect,    //                        .chipselect
		input  wire        onchip_memory2_0_s1_write,         //                        .write
		output wire [7:0]  onchip_memory2_0_s1_readdata,      //                        .readdata
		input  wire [7:0]  onchip_memory2_0_s1_writedata      //                        .writedata
	);

	background_data_onchip_memory2_0 onchip_memory2_0 (
		.clk         (onchip_memory2_0_clk1_clk),         //   clk1.clk
		.address     (onchip_memory2_0_s1_address),       //     s1.address
		.debugaccess (onchip_memory2_0_s1_debugaccess),   //       .debugaccess
		.clken       (onchip_memory2_0_s1_clken),         //       .clken
		.chipselect  (onchip_memory2_0_s1_chipselect),    //       .chipselect
		.write       (onchip_memory2_0_s1_write),         //       .write
		.readdata    (onchip_memory2_0_s1_readdata),      //       .readdata
		.writedata   (onchip_memory2_0_s1_writedata),     //       .writedata
		.reset       (onchip_memory2_0_reset1_reset),     // reset1.reset
		.reset_req   (onchip_memory2_0_reset1_reset_req), //       .reset_req
		.freeze      (1'b0)                               // (terminated)
	);

endmodule
