// audio_system.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module audio_system (
		input  wire        audio_0_external_interface_ADCDAT,                           //                      audio_0_external_interface.ADCDAT
		input  wire        audio_0_external_interface_ADCLRCK,                          //                                                .ADCLRCK
		input  wire        audio_0_external_interface_BCLK,                             //                                                .BCLK
		output wire        audio_0_external_interface_DACDAT,                           //                                                .DACDAT
		input  wire        audio_0_external_interface_DACLRCK,                          //                                                .DACLRCK
		input  wire [1:0]  audio_and_video_config_0_avalon_av_config_slave_address,     // audio_and_video_config_0_avalon_av_config_slave.address
		input  wire [3:0]  audio_and_video_config_0_avalon_av_config_slave_byteenable,  //                                                .byteenable
		input  wire        audio_and_video_config_0_avalon_av_config_slave_read,        //                                                .read
		input  wire        audio_and_video_config_0_avalon_av_config_slave_write,       //                                                .write
		input  wire [31:0] audio_and_video_config_0_avalon_av_config_slave_writedata,   //                                                .writedata
		output wire [31:0] audio_and_video_config_0_avalon_av_config_slave_readdata,    //                                                .readdata
		output wire        audio_and_video_config_0_avalon_av_config_slave_waitrequest, //                                                .waitrequest
		inout  wire        audio_and_video_config_0_external_interface_SDAT,            //     audio_and_video_config_0_external_interface.SDAT
		output wire        audio_and_video_config_0_external_interface_SCLK,            //                                                .SCLK
		output wire        audio_final_fifo_almost_empty_data,                          //                   audio_final_fifo_almost_empty.data
		output wire        audio_final_fifo_almost_full_data,                           //                    audio_final_fifo_almost_full.data
		input  wire [15:0] audio_final_fifo_in_data,                                    //                             audio_final_fifo_in.data
		input  wire        audio_final_fifo_in_valid,                                   //                                                .valid
		output wire        audio_final_fifo_in_ready,                                   //                                                .ready
		output wire [15:0] audio_final_fifo_out_data,                                   //                            audio_final_fifo_out.data
		output wire        audio_final_fifo_out_valid,                                  //                                                .valid
		input  wire        audio_final_fifo_out_ready,                                  //                                                .ready
		output wire        audio_pll_0_audio_clk_clk,                                   //                           audio_pll_0_audio_clk.clk
		output wire        audio_sc_fifo_almost_empty_data,                             //                      audio_sc_fifo_almost_empty.data
		output wire        audio_sc_fifo_almost_full_data,                              //                       audio_sc_fifo_almost_full.data
		output wire [15:0] audio_sc_fifo_out_data,                                      //                               audio_sc_fifo_out.data
		output wire        audio_sc_fifo_out_valid,                                     //                                                .valid
		input  wire        audio_sc_fifo_out_ready,                                     //                                                .ready
		input  wire        clk_clk,                                                     //                                             clk.clk
		input  wire        reset_reset_n                                                //                                           reset.reset_n
	);

	wire         audio_0_avalon_left_channel_source_valid;  // audio_0:from_adc_left_channel_valid -> audio_sc_fifo:in_valid
	wire  [15:0] audio_0_avalon_left_channel_source_data;   // audio_0:from_adc_left_channel_data -> audio_sc_fifo:in_data
	wire         audio_0_avalon_left_channel_source_ready;  // audio_sc_fifo:in_ready -> audio_0:from_adc_left_channel_ready
	wire         audio_0_avalon_right_channel_source_valid; // audio_0:from_adc_right_channel_valid -> audio_0:to_dac_right_channel_valid
	wire  [15:0] audio_0_avalon_right_channel_source_data;  // audio_0:from_adc_right_channel_data -> audio_0:to_dac_right_channel_data
	wire         audio_0_avalon_right_channel_source_ready; // audio_0:to_dac_right_channel_ready -> audio_0:from_adc_right_channel_ready
	wire         rst_controller_reset_out_reset;            // rst_controller:reset_out -> [audio_0:reset, audio_and_video_config_0:reset, audio_sc_fifo:reset]
	wire         audio_pll_0_reset_source_reset;            // audio_pll_0:reset_source_reset -> rst_controller:reset_in0
	wire         rst_controller_001_reset_out_reset;        // rst_controller_001:reset_out -> audio_final_fifo:reset

	audio_system_audio_0 audio_0 (
		.clk                          (clk_clk),                                   //                         clk.clk
		.reset                        (rst_controller_reset_out_reset),            //                       reset.reset
		.from_adc_left_channel_ready  (audio_0_avalon_left_channel_source_ready),  //  avalon_left_channel_source.ready
		.from_adc_left_channel_data   (audio_0_avalon_left_channel_source_data),   //                            .data
		.from_adc_left_channel_valid  (audio_0_avalon_left_channel_source_valid),  //                            .valid
		.from_adc_right_channel_ready (audio_0_avalon_right_channel_source_ready), // avalon_right_channel_source.ready
		.from_adc_right_channel_data  (audio_0_avalon_right_channel_source_data),  //                            .data
		.from_adc_right_channel_valid (audio_0_avalon_right_channel_source_valid), //                            .valid
		.to_dac_left_channel_data     (),                                          //    avalon_left_channel_sink.data
		.to_dac_left_channel_valid    (),                                          //                            .valid
		.to_dac_left_channel_ready    (),                                          //                            .ready
		.to_dac_right_channel_data    (audio_0_avalon_right_channel_source_data),  //   avalon_right_channel_sink.data
		.to_dac_right_channel_valid   (audio_0_avalon_right_channel_source_valid), //                            .valid
		.to_dac_right_channel_ready   (audio_0_avalon_right_channel_source_ready), //                            .ready
		.AUD_ADCDAT                   (audio_0_external_interface_ADCDAT),         //          external_interface.export
		.AUD_ADCLRCK                  (audio_0_external_interface_ADCLRCK),        //                            .export
		.AUD_BCLK                     (audio_0_external_interface_BCLK),           //                            .export
		.AUD_DACDAT                   (audio_0_external_interface_DACDAT),         //                            .export
		.AUD_DACLRCK                  (audio_0_external_interface_DACLRCK)         //                            .export
	);

	audio_system_audio_and_video_config_0 audio_and_video_config_0 (
		.clk         (clk_clk),                                                     //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                              //                  reset.reset
		.address     (audio_and_video_config_0_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (audio_and_video_config_0_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (audio_and_video_config_0_avalon_av_config_slave_read),        //                       .read
		.write       (audio_and_video_config_0_avalon_av_config_slave_write),       //                       .write
		.writedata   (audio_and_video_config_0_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (audio_and_video_config_0_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (audio_and_video_config_0_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (audio_and_video_config_0_external_interface_SDAT),            //     external_interface.export
		.I2C_SCLK    (audio_and_video_config_0_external_interface_SCLK)             //                       .export
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (2),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (65536),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (1),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (1),
		.USE_ALMOST_EMPTY_IF (1)
	) audio_final_fifo (
		.clk               (clk_clk),                            //          clk.clk
		.reset             (rst_controller_001_reset_out_reset), //    clk_reset.reset
		.csr_address       (),                                   //          csr.address
		.csr_read          (),                                   //             .read
		.csr_write         (),                                   //             .write
		.csr_readdata      (),                                   //             .readdata
		.csr_writedata     (),                                   //             .writedata
		.almost_full_data  (audio_final_fifo_almost_full_data),  //  almost_full.data
		.almost_empty_data (audio_final_fifo_almost_empty_data), // almost_empty.data
		.in_data           (audio_final_fifo_in_data),           //           in.data
		.in_valid          (audio_final_fifo_in_valid),          //             .valid
		.in_ready          (audio_final_fifo_in_ready),          //             .ready
		.out_data          (audio_final_fifo_out_data),          //          out.data
		.out_valid         (audio_final_fifo_out_valid),         //             .valid
		.out_ready         (audio_final_fifo_out_ready),         //             .ready
		.in_startofpacket  (1'b0),                               //  (terminated)
		.in_endofpacket    (1'b0),                               //  (terminated)
		.out_startofpacket (),                                   //  (terminated)
		.out_endofpacket   (),                                   //  (terminated)
		.in_empty          (1'b0),                               //  (terminated)
		.out_empty         (),                                   //  (terminated)
		.in_error          (1'b0),                               //  (terminated)
		.out_error         (),                                   //  (terminated)
		.in_channel        (1'b0),                               //  (terminated)
		.out_channel       ()                                    //  (terminated)
	);

	audio_system_audio_pll_0 audio_pll_0 (
		.ref_clk_clk        (clk_clk),                        //      ref_clk.clk
		.ref_reset_reset    (~reset_reset_n),                 //    ref_reset.reset
		.audio_clk_clk      (audio_pll_0_audio_clk_clk),      //    audio_clk.clk
		.reset_source_reset (audio_pll_0_reset_source_reset)  // reset_source.reset
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (2),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (1),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (1),
		.USE_ALMOST_EMPTY_IF (1)
	) audio_sc_fifo (
		.clk               (clk_clk),                                  //          clk.clk
		.reset             (rst_controller_reset_out_reset),           //    clk_reset.reset
		.csr_address       (),                                         //          csr.address
		.csr_read          (),                                         //             .read
		.csr_write         (),                                         //             .write
		.csr_readdata      (),                                         //             .readdata
		.csr_writedata     (),                                         //             .writedata
		.almost_full_data  (audio_sc_fifo_almost_full_data),           //  almost_full.data
		.almost_empty_data (audio_sc_fifo_almost_empty_data),          // almost_empty.data
		.in_data           (audio_0_avalon_left_channel_source_data),  //           in.data
		.in_valid          (audio_0_avalon_left_channel_source_valid), //             .valid
		.in_ready          (audio_0_avalon_left_channel_source_ready), //             .ready
		.out_data          (audio_sc_fifo_out_data),                   //          out.data
		.out_valid         (audio_sc_fifo_out_valid),                  //             .valid
		.out_ready         (audio_sc_fifo_out_ready),                  //             .ready
		.in_startofpacket  (1'b0),                                     //  (terminated)
		.in_endofpacket    (1'b0),                                     //  (terminated)
		.out_startofpacket (),                                         //  (terminated)
		.out_endofpacket   (),                                         //  (terminated)
		.in_empty          (1'b0),                                     //  (terminated)
		.out_empty         (),                                         //  (terminated)
		.in_error          (1'b0),                                     //  (terminated)
		.out_error         (),                                         //  (terminated)
		.in_channel        (1'b0),                                     //  (terminated)
		.out_channel       ()                                          //  (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (audio_pll_0_reset_source_reset), // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
